`timescale 1ns / 1ps


module ROT_Cordic
#(parameter M=32,N=5)
(input signed [M-1:0] x_in,
 input signed [M-1:0] y_in,
 input signed [M-1:0] z_in,
 input [1:0] mode,
 input clk,
 input rst,
 output signed [M-1:0] xf,
 output signed [M-1:0] yf,
 output signed [M-1:0] zf);
 
 genvar j;
 
 wire signed [M-1:0] x [0:M];
 wire signed [M-1:0] y [0:M];
 wire signed [M-1:0] z [0:M];
 
// localparam signed [M-1:0] pi_2=32'b00110010010000111111011010101001;
// localparam signed [M-1:0] minus_pi_2 = 32'b11001101101111000000100101010111;
 
 wire signed [31:0] atanj [0:M-1];

assign atanj[0]  = (mode[1]) ? 32'b00010001100100111110101001111011 : 32'b00011001000111111011010101000100;
assign atanj[1]  = (mode[1]) ? 32'b00001000001011000101011101111101 : 32'b00001110110101100011100101111001;
assign atanj[2]  = (mode[1]) ? 32'b00000100000001010110001001000111 : 32'b00000111110101101101101110110011;
assign atanj[3]  = (mode[1]) ? 32'b00000010000000001010101100010001 : 32'b00000011111101011010111110011100;
assign atanj[4]  = (mode[1]) ? 32'b00000001000000000001010101011001 : 32'b00000001111111101010111001010010;
assign atanj[5]  = (mode[1]) ? 32'b00000000100000000000001010101011 : 32'b00000000111111111101010111011000;
assign atanj[6]  = (mode[1]) ? 32'b00000000010000000000000001010101 : 32'b00000000011111111111101010111011;
assign atanj[7]  = (mode[1]) ? 32'b00000000001000000000000000001011 : 32'b00000000001111111111111101010111;
assign atanj[8]  = (mode[1]) ? 32'b00000000000100000000000000000001 : 32'b00000000000111111111111111101011;
assign atanj[9]  = (mode[1]) ? 32'b00000000000010000000000000000000 : 32'b00000000000011111111111111111101;
assign atanj[10] = (mode[1]) ? 32'b00000000000001000000000000000000 : 32'b00000000000001111111111111111111;
assign atanj[11] = (mode[1]) ? 32'b00000000000000100000000000000000 : 32'b00000000000000111111111111111111;
assign atanj[12] = (mode[1]) ? 32'b00000000000000010000000000000000 : 32'b00000000000000011111111111111111;
assign atanj[13] = (mode[1]) ? 32'b00000000000000001000000000000000 : 32'b00000000000000001111111111111111;
assign atanj[14] = (mode[1]) ? 32'b00000000000000000100000000000000 : 32'b00000000000000000111111111111111;
assign atanj[15] = (mode[1]) ? 32'b00000000000000000010000000000000 : 32'b00000000000000000011111111111111;
assign atanj[16] = (mode[1]) ? 32'b00000000000000000001000000000000 : 32'b00000000000000000001111111111111;
assign atanj[17] = (mode[1]) ? 32'b00000000000000000000100000000000 : 32'b00000000000000000000111111111111;
assign atanj[18] = (mode[1]) ? 32'b00000000000000000000010000000000 : 32'b00000000000000000000011111111111;
assign atanj[19] = (mode[1]) ? 32'b00000000000000000000001000000000 : 32'b00000000000000000000001111111111;
assign atanj[20] = (mode[1]) ? 32'b00000000000000000000000100000000 : 32'b00000000000000000000000111111111;
assign atanj[21] = (mode[1]) ? 32'b00000000000000000000000010000000 : 32'b00000000000000000000000011111111;
assign atanj[22] = (mode[1]) ? 32'b00000000000000000000000001000000 : 32'b00000000000000000000000001111111;
assign atanj[23] = (mode[1]) ? 32'b00000000000000000000000000100000 : 32'b00000000000000000000000000111111;
assign atanj[24] = (mode[1]) ? 32'b00000000000000000000000000010000 : 32'b00000000000000000000000000011111;
assign atanj[25] = (mode[1]) ? 32'b00000000000000000000000000001000 : 32'b00000000000000000000000000001111;
assign atanj[26] = (mode[1]) ? 32'b00000000000000000000000000000100 : 32'b00000000000000000000000000000111;
assign atanj[27] = (mode[1]) ? 32'b00000000000000000000000000000010 : 32'b00000000000000000000000000000011;
assign atanj[28] = (mode[1]) ? 32'b00000000000000000000000000000001 : 32'b00000000000000000000000000000001;
assign atanj[29] = (mode[1]) ? 32'b00000000000000000000000000000000 : 32'b00000000000000000000000000000000;
assign atanj[30] = (mode[1]) ? 32'b00000000000000000000000000000000 : 32'b00000000000000000000000000000000;
assign atanj[31] = (mode[1]) ? 32'b00000000000000000000000000000000 : 32'b00000000000000000000000000000000;

pre_stage m1(x_in,y_in,z_in,mode,clk,x[0],y[0],z[0]);

assign xf = x[M];
assign yf = y[M];
assign zf = z[M];
    
 generate
 for( j=0; j<M; j=j+1)
 begin
 Cordic_stage c1 (x[j],y[j],z[j],mode,rst,atanj[j],j,clk,x[j+1],y[j+1],z[j+1]);
 end 
 endgenerate
endmodule
